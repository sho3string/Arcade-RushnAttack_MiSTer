//----------------------------------
//  Dual-Port RAM for VIDEO
//----------------------------------
// Copyright (c) 2013,19 MiSTer-X

module VRAM4096
(
	input					cl,
	input	 [11:0]		ad,
	input					en,
	input					wr,
	input   [7:0]		id,
	output reg [7:0]	od,

	input					clv,
	input  [11:0]		adv,
	output reg [7:0]	odv
);

reg [7:0] core [0:4095];

always @( posedge cl ) begin
	if (en) begin
		if (wr) core[ad] <= id;
		else od <= core[ad];
	end
end

always @( posedge clv ) begin
	odv <= core[adv];
end

endmodule

module VRAM2048
(
	input					cl,
	input	 [10:0]		ad,
	input					en,
	input					wr,
	input   [7:0]		id,
	output reg [7:0]	od,

	input					clv,
	input  [10:0]		adv,
	output reg [7:0]	odv
);

reg [7:0] core [0:2047];

always @( posedge cl ) begin
	if (en) begin
		if (wr) core[ad] <= id;
		else od <= core[ad];
	end
end

always @( posedge clv ) begin
	odv <= core[adv];
end

endmodule

module VRAM32
(
	input					cl,
	input	  [4:0]		ad,
	input					en,
	input					wr,
	input   [7:0]		id,
	output reg [7:0]	od,

	input					clv,
	input   [4:0]		adv,
	output reg [7:0]	odv
);

reg [7:0] core [0:31];

always @( posedge cl ) begin
	if (en) begin
		if (wr) core[ad] <= id;
		else od <= core[ad];
	end
end

always @( posedge clv ) begin
	odv <= core[adv];
end

endmodule


module LineBuf
(
	input				WCL,
	input				WEN,
	input	 [9:0]	WAD,
	input  [3:0]	WDT,

	input				RCL,
	input				RWE,
	input  [9:0]	RAD,
	output reg [3:0]	RDT
);

wire [3:0] dum;

reg [10:0] ram[0:1023];

always @(posedge RCL) begin
	if(RWE) begin
		ram[RAD] <= 0;
		RDT <= 0;
	end
	else begin
		RDT <= ram[RAD];
	end
end

always @(posedge WCL) begin
	if(WEN) begin
		ram[WAD] <= WDT;
	end
end

/*
DPRAM1024_4 ramcore
(
	WAD, RAD,
	WCL, RCL,
	WDT, 4'h0,
	WEN, RWE,
	dum, RDT
);*/

endmodule

